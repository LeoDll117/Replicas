----------------------------------------------------------------------------------
--Ejercicio contador asc-desc carga paralelo pagina 64
--Leonardo Peralta
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_arith.all;
use IEEE.STD_LOGIC_SIGNED.ALL;

entity contador5 is
    Port ( clk, LD, UP : in  STD_LOGIC;
           D : in  STD_LOGIC_VECTOR (2 downto 0);
           Q : inout  STD_LOGIC_VECTOR (2 downto 0));
end contador5;

architecture modulo of contador5 is
begin
	process(clk, LD, D, UP) 
		begin
			if(clk' event and clk='1')then
				if(LD ='0')then
					Q<=D;
				elsif UP ='1' then
					Q <= Q+1;
				else
					Q<=Q-1;
				end if;
			end if;
		end process;
	end modulo; 
				
	
